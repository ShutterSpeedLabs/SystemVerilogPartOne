class second;

  constraint data_c_s {data_s > 10; data_s < 20;}
  rand int data_s;
  
endclass
