class first;
  
  rand int data;
  
  constraint data_c {data < 10; data > 0;}
 
endclass
