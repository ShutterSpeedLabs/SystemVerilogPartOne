class transaction;
  
  bit [7:0] data;
  
endclass
