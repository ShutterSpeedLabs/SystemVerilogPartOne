class generator;
  
  rand bit [3:0] a, b; ////////////rand or randc 
  
endclass