class transaction;
  
    rand bit [7:0] a;
    rand bit [7:0] b;
    rand bit wr;
 
endclass
