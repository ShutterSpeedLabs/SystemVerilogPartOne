class first;
  
  constraint data_c_f { data_f > 0; data_f < 10;}
  rand int data_f;
   
endclass
