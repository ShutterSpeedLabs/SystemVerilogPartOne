class second;
  
  rand int data;
  
  constraint data_c {data > 10; data < 20;}
  
endclass
